module main

fn main() {
	println(Buffer.from_int64learray([i64(-128)]))
}